module FPMUL (
  input wire CLK,
  input wire RST_N,
  input wire [7:0] A,
  input wire [7:0] B,
  input wire START,
  output reg [7:0] Y,
  output reg signed [4:0] E,
  output reg DONE
);

  // Write your code here

endmodule
